module Hazard_Unit();
endmodule