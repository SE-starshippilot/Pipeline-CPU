module Flush();

endmodule